/* 
	Description : Component convolution_1_1 which perform the 1*1 convolution needed for inverted residual block and 1*1 convolution layer
	Author : 	  Guillaume Gheysen
*/ 

/* 
	###################################################################################################################################
	# import 																																								 #
   ###################################################################################################################################
*/
import dma_pkg::*;
import ram_pkg::*;
/* 
	###################################################################################################################################
	# module definition 																																					 #
   ###################################################################################################################################
*/
module Convolution_1_1(input logic clk, rst, start,
							  input logic signed [PX_W - 1:0] fmi_data,
							  input logic signed [WG_W -1:0] kex_data,
							  input logic [$clog2(Npar) - 1:0] kex_pos,
							  input logic [10:0] Nif,
							  output logic [$clog2(FMI_N_ELEM)-1:0] fmi_addr,
							  output logic [$clog2(KEX_N_ELEM)-1:0] kex_addr,
							  output logic [$clog2(FMINT_N_ELEM)-1:0] fmint_addr,
							  output logic finish, write,
							  output logic signed [PX_W - 1:0] res
							 );
	
	/* 
		###################################################################################################################################
		# internal signals																																					 #
		###################################################################################################################################
	*/
	// States
	typedef enum logic [2:0] {IDLE,             
									  FINISHED,					// State telling the DMA has finished its transaction
									  LOAD_DATA,
									  FINISHED_LOAD,
									  COMPUTATION,
									  WRITE
									  } statetype;
	statetype state, state_n; // Variables containing the state
	
	// Registers
	logic signed [PX_W - 1:0]  px  [Npar-1 : 0];
	logic signed [WG_W - 1:0]  wg  [Nnp-1 : 0];
	logic [$clog2(Npar) - 1:0] pos [Nnp-1 : 0];
	logic [7:0] x_fmi, y_fmi;
	logic [10:0] f_fmi, f_fmint, tf_fmi;
	logic [10:0] np_kex;
	logic [$clog2(FMI_N_ELEM)-1:0] fmi_addr_ref;
	logic [$clog2(KEX_N_ELEM)-1:0] f_kex_mem;
	logic load_px, load_wg;
	logic signed [PX_W - 1:0] sum;
	// Next value for registers 
	logic [7:0] x_fmi_n, y_fmi_n;
	logic [10:0] f_fmi_n, f_fmint_n, tf_fmi_n;
	logic [$clog2(FMI_N_ELEM)-1:0] fmi_addr_n, fmi_addr_ref_n;
	logic [$clog2(FMINT_N_ELEM)-1:0] fmint_addr_n;
	logic [10:0] np_kex_n;
	logic [$clog2(KEX_N_ELEM)-1:0] kex_addr_n, f_kex_mem_n;
	logic load_px_n, load_wg_n;
	logic signed [PX_W - 1:0] sum_n; 
	 
	/* 
		###################################################################################################################################
		# Modules instatiation																																					 #
		###################################################################################################################################
	*/
	SHIFT_REGISTER_PX reg_px(.clk(clk), .load(load_px), .data(fmi_data), .pixels(px));
	SHIFT_REGISTER_WG reg_wg(.clk(clk), .load(load_wg), .data(kex_data), .weights(wg));
	SHIFT_REGISTER_POS reg_pos(.clk(clk), .load(load_wg), .data(kex_pos), .pos(pos));
	
	RELU6 activation(.in(sum), .out(res));
	
	/* 
		###################################################################################################################################
		# Sequential logic																																					 #
		###################################################################################################################################
	*/
	always_ff @(posedge clk, posedge rst) begin
		if(rst) begin
			state <= IDLE;
			x_fmi <= '0; y_fmi <= '0;
			f_fmi <= '0; f_fmint <= '0; tf_fmi <= '0;
			fmint_addr <= '0; fmi_addr <= '0; fmi_addr_ref <= '0;
			np_kex <= '0;
			kex_addr <= '0; f_kex_mem <= '0;
			load_px <= '0; load_wg <= '0;
			sum <= '0;
		end
		else begin
			state <= state_n;
			x_fmi <= x_fmi_n; y_fmi <= y_fmi_n;
			f_fmi <= f_fmi_n; f_fmint <= f_fmint_n; tf_fmi <= tf_fmi_n;
			fmint_addr <= fmint_addr_n; 
			fmi_addr <= fmi_addr_n; 
			fmi_addr_ref <= fmi_addr_ref_n;
			np_kex <= np_kex_n;
			kex_addr <= kex_addr_n;
			f_kex_mem <= f_kex_mem_n;
			load_px <= load_px_n; 
			load_wg <= load_wg_n;
			sum <= sum_n;
		end
	end
	
	/* 
		###################################################################################################################################
		# Combinational logic																																				 #
		###################################################################################################################################
	*/
	assign finish = state == FINISHED;
	assign write = state == WRITE;
	
	always_comb begin
		state_n = state;
		x_fmi_n = x_fmi; y_fmi_n = y_fmi;
		f_fmi_n = f_fmi; f_fmint_n = f_fmint; tf_fmi_n = tf_fmi;
		fmint_addr_n = fmint_addr; 
		fmi_addr_n = fmi_addr; 
		fmi_addr_ref_n = fmi_addr_ref;
		np_kex_n = np_kex;
		kex_addr_n = kex_addr; f_kex_mem_n = f_kex_mem;
		load_px_n = load_px; load_wg_n = load_wg;
		sum_n = sum;
		case(state) 
			// IDLE state - when no computation is occuring
			IDLE: begin
				if(start) begin
					state_n = LOAD_DATA;
					// FMI variables
					x_fmi_n = 1; y_fmi_n = 1; f_fmint_n = 1; fmint_addr_n = '0; // Output pixels variables & address
					f_fmi_n = 1; tf_fmi_n = 1; fmi_addr_n = '0; fmi_addr_ref_n = '0;// FMI variables
					// KEX variables
					np_kex_n = 1;
					kex_addr_n = '0; f_kex_mem_n = '0;// 
					// Sum
					sum_n = '0;
				end
			end
			
			// IDLE state - when the component has finished its computation
		   FINISHED: begin
				state_n = IDLE;
			end
			
		   LOAD_DATA: begin
				if (tf_fmi == Npar - 1|| f_fmi == Nif - 1 ) begin
					state_n = FINISHED_LOAD;
					load_px_n = '1;
					f_fmi_n = f_fmi + 11'b1;
					tf_fmi_n = tf_fmi + 11'b1;
				end
				else begin
					load_px_n = 'b1;
					f_fmi_n = f_fmi + load_px;
					tf_fmi_n = tf_fmi + load_px;
					fmi_addr_n = fmi_addr + FMI_N_CHAN[$clog2(FMI_N_ELEM)-1:0];
				end
				
				if (np_kex == Nnp) begin
					if(np_kex == 1) begin
						load_wg_n = 1;
					end
					else begin
						load_wg_n = 0;
					end
				end
				else if (np_kex == Nnp - 1) begin
					load_wg_n = '1; 
					np_kex_n = np_kex + load_wg;
					kex_addr_n = kex_addr + {{$clog2(KEX_N_ELEM) - 1{1'b0}}, ~load_wg}; 
				end
				else begin
					load_wg_n = 1;
					np_kex_n = np_kex + load_wg;
					kex_addr_n = kex_addr + {{$clog2(KEX_N_ELEM) - 1{1'b0}}, 1'b1};
				end
			end
			
			FINISHED_LOAD: begin
				state_n = COMPUTATION;
				load_px_n = '0;
				load_wg_n = '0; 
			end
		
		   COMPUTATION: begin
				for(int i = 0; i < Nnp ; i=i+1) begin
					// Intermediate values
					logic signed [PX_W - 1 : 0] cur_val;
					logic signed [WG_W - 1 : 0] cur_wg;
					logic signed [$clog2(Npar):0] cur_pos;
					logic signed [(2*PX_W) - 1 : 0] int_res;
					logic signed [PX_W - 1 : 0] trunc_res;
					logic signed [PX_W - 1 : 0] round_res;
					// COmputation
					cur_pos[$clog2(Npar)-1:0] = pos[i][$clog2(Npar) -1 :0];
					cur_val = px[cur_pos[$clog2(Npar)-1:0]][PX_W - 1 : 0];
					cur_wg = wg[i][WG_W - 1:0];
					int_res = cur_val * cur_wg;
					trunc_res = int_res[(2*PX_W) - 4 - 1: PX_W - 4];
					round_res = int_res[(2*PX_W) - 4 - 1];
					sum_n = sum_n + trunc_res + round_res; 
				end
				if(f_fmi == Nif) begin
					state_n = WRITE;
				end
				else begin
					state_n = LOAD_DATA;
					f_fmi_n = f_fmi + 11'b1;
					tf_fmi_n = 1; 
					fmi_addr_n = fmi_addr + FMI_N_CHAN[$clog2(FMI_N_ELEM)-1:0]; // We change the Par (next channel)
					np_kex_n = 1; kex_addr_n = kex_addr + '1; // We change the group (next weight)
				end
			end
			
		   WRITE: begin
				fmint_addr_n = fmint_addr + {{$clog2(FMINT_N_ELEM) - 1{1'b0}}, 1'b1};
				sum_n = '0;
				f_fmi_n = 1;
				if (x_fmi == Tix) begin // Change column
					x_fmi_n = 1;
					if (y_fmi == Tiy) begin // Change row
						y_fmi_n = 1; fmi_addr_n = '0; fmi_addr_ref_n = '0;
						if (f_fmint == Npar) begin
							state_n = FINISHED;
						end
						else begin // Kernel change
							state_n = LOAD_DATA;
							f_fmint_n = f_fmint + 11'b1;
							kex_addr_n = kex_addr + {{$clog2(KEX_N_ELEM) - 1{1'b0}}, 1'b1};
							f_kex_mem_n = kex_addr + {{$clog2(KEX_N_ELEM) - 1{1'b0}}, 1'b1};
							np_kex_n = 1;
						end
					end
					else begin // Spatial change
						state_n = LOAD_DATA;
						y_fmi_n = y_fmi + 8'b1;
						tf_fmi_n = 1; 	
						fmi_addr_n = fmi_addr_ref + {{$clog2(FMI_N_ELEM) - 1{1'b0}}, 1'b1};
						fmi_addr_ref_n = fmi_addr_ref + {{$clog2(FMI_N_ELEM) - 1{1'b0}}, 1'b1};
						kex_addr_n = f_kex_mem;
						np_kex_n = 1;
					end
				end
				else begin // Spatial change
					state_n = LOAD_DATA;
					x_fmi_n = x_fmi + 8'b1;
					tf_fmi_n = 1; 
					fmi_addr_n = fmi_addr_ref + {{$clog2(FMI_N_ELEM) - 1{1'b0}}, 1'b1};
					fmi_addr_ref_n = fmi_addr_ref + {{$clog2(FMI_N_ELEM) - 1{1'b0}}, 1'b1};
					kex_addr_n = f_kex_mem;
					np_kex_n = 1;
				end
			end
		endcase
	end
endmodule
/* 
	###################################################################################################################################
	# Additional modules																																				 #
	###################################################################################################################################
*/
module SHIFT_REGISTER_PX(
								 input logic clk, load,
								 input logic signed[PX_W - 1:0] data,
								 output logic signed [PX_W - 1:0] pixels [Npar-1 : 0]
								);
	always_ff @(posedge clk) begin
		if (load) begin
		pixels [Npar-1] <= data;
		for (int i=0 ; i < Npar -1; i=i+1) begin
			pixels[i] <= pixels[i+1];
		end
		end
	end
endmodule

module SHIFT_REGISTER_WG(
								 input logic clk, load,
								 input logic signed [WG_W  - 1:0] data,
								 output logic signed [WG_W  - 1:0] weights [Nnp-1 : 0]
								);
	always_ff @(posedge clk) begin
		if (load) begin
		weights [Nnp-1] <= data;
		for (int i=0 ; i < Nnp-1; i=i+1) begin
			weights[i] <= weights[i+1];
		end
		end
	end
endmodule

module SHIFT_REGISTER_POS(
								 input logic clk, load,
								 input logic [$clog2(Npar) - 1:0] data,
								 output logic [$clog2(Npar) - 1:0] pos [Nnp-1 : 0]
								);
	always_ff @(posedge clk) begin
		if (load) begin
			pos [Nnp-1] <= data;
				for (int i=0 ; i < Nnp-1; i=i+1) begin
					pos[i] <= pos[i+1];
				end
			end
	end
endmodule

module RELU6(
				 input logic signed [PX_W - 1:0] in,
				 output logic signed [PX_W - 1:0] out);
	logic [PX_W -1 : 0] val = (4'b0110) << (PX_W - 4 - 1);
	assign out = in[PX_W - 1] ? '0 : ( (in[PX_W - 1:PX_W - 4 -1] == 4'b0110) ? val : in);
endmodule
