/* 
	Description : RAM component, containing the tile of the kernels of DW convolution
	Author : 	  Guillaume Gheysen
*/
 
/* 
	###################################################################################################################################
	# import 																																								 #
   ###################################################################################################################################
*/
import irb_pkg::*;
/* 
	###################################################################################################################################
	# module definition 																																					 #
   ###################################################################################################################################
*/
module RAM_KDW(
						input logic  clk,									  // Clock
						input logic  [$clog2(KDW_N_ELEM+1)-1:0] addr, // Ram address to read/write data
						input logic  [WG_W -1:0] data,				  // if write is enabled, data to write at address addr
						input logic  write,								  // if enabled, write data
						output logic [WG_W-1:0] res					  // Data
					);
	/* 
		################################################################################################################################
		# RAM 																																			            	 #
		################################################################################################################################
	*/
	logic [WG_W-1:0] mem [0:KDW_N_ELEM-1];
	/* 
		################################################################################################################################
		# Sequential logic																																				 #
		################################################################################################################################
	*/
	always_ff @(posedge clk) begin
		if (write) begin
			mem[addr] <= data;
			res <= data;
		end 
		else res <= mem[addr];
	end
endmodule
