
module RAM(
	input logic clk,
	input logic [2:0] addr,
	input logic [15:0] data,
	input logic write,
	output logic [15:0] res);
	
	logic [15:0] mem [7:0];

	always_ff @(posedge clk) begin
	if (write) begin
		mem[addr] <= data;
		res <= data;
	end 
	else res <= mem[addr];
	end
endmodule
