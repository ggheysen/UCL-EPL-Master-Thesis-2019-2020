/* 
	Description : RAM component, containing the tile of FM output
	Author : 	  Guillaume Gheysen
*/
 
/* 
	###################################################################################################################################
	# import 																																								 #
   ###################################################################################################################################
*/
import irb_pkg::*;
/* 
	###################################################################################################################################
	# module definition 																																					 #
   ###################################################################################################################################
*/
module RAM_FMO(
						input logic  clk, 								  // Clock
						input logic  [$clog2(FMO_N_ELEM)-1:0] addr, // Ram address to read/write data
						input logic  [PX_W-1:0] data,					  // if write is enabled, data to write at address addr
						input logic  write,								  // if enabled, write data
						output logic [PX_W-1:0] res					  // Data
					);
	/* 
		################################################################################################################################
		# RAM 																																			            	 #
		################################################################################################################################
	*/
	logic [PX_W-1:0] mem [FMO_N_ELEM-1:0];
	/* 
		################################################################################################################################
		# Sequential logic																																				 #
		################################################################################################################################
	*/
	always_ff @(posedge clk) begin
		if (write) begin
			mem[addr] <= data;
			res <= data;
		end 
		else res <= mem[addr];
	end
endmodule
