/* 
	Description : RAM component, containing the tile of FM of intermediate result
	Author : 	  Guillaume Gheysen
*/
 
/* 
	###################################################################################################################################
	# import 																																								 #
   ###################################################################################################################################
*/
import irb_pkg::*;

/* 
	###################################################################################################################################
	# module definition 																																					 #
   ###################################################################################################################################
*/
module RAM_FMINT(
						input logic  clk, 									 // Clock
						input logic  [$clog2(FMINT_N_ELEM)-1:0] addr, // Ram address to read/write data
						input logic  [PX_W-1:0] data,						 // if write is enabled, data to write at address addr
						input logic  write,									 // if enabled, write data
						output logic [PX_W-1:0] res						 // Data
					);

	/* 
		################################################################################################################################
		# RAM 																																			            	 #
		################################################################################################################################
	*/	
	logic [PX_W-1:0] mem [FMINT_N_ELEM-1:0];
	/* 
		################################################################################################################################
		# Sequential logic																																				 #
		################################################################################################################################
	*/
	always_ff @(posedge clk) begin
		if (write) begin
			mem[addr] <= data;
			res <= data;
		end 
		else res <= mem[addr];
	end
endmodule
